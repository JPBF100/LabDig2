module sonar (
 input clock,
 input reset,
 input ligar,
 input echo,
 output trigger,
 output pwm,
 output saida_serial,
 output fim_posição
); 


endmodule