module sonar (
 input wire clock,
 input wire reset,
 input wire ligar,
 input wire echo,
 output wire trigger,
 output wire pwm,
 output wire saida_serial,
 output wire fim_posição
); 

endmodule